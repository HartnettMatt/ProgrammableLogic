// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// Created on Sun Oct 29 21:38:51 2023

// synthesis message_off 10175

`timescale 1ns/1ns

module HW3Q6 (
    reset,clock,A,B,C,D,PBGNT,MACK,CONT,
    PBREQ,CMREQ,CE,CNTLD);

    input reset;
    input clock;
    input A;
    input B;
    input C;
    input D;
    input PBGNT;
    input MACK;
    input CONT;
    tri0 reset;
    tri0 A;
    tri0 B;
    tri0 C;
    tri0 D;
    tri0 PBGNT;
    tri0 MACK;
    tri0 CONT;
    output PBREQ;
    output CMREQ;
    output CE;
    output CNTLD;
    reg PBREQ;
    reg CMREQ;
    reg CE;
    reg CNTLD;
    reg [5:0] fstate;
    reg [5:0] reg_fstate;
    parameter state0=0,state3=1,state1=2,state2=3,state4=4,state5=5;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or A or B or C or D or PBGNT or MACK or CONT)
    begin
        if (reset) begin
            reg_fstate <= state0;
            PBREQ <= 1'b0;
            CMREQ <= 1'b0;
            CE <= 1'b0;
            CNTLD <= 1'b0;
        end
        else begin
            PBREQ <= 1'b0;
            CMREQ <= 1'b0;
            CE <= 1'b0;
            CNTLD <= 1'b0;
            case (fstate)
                state0: begin
                    if ((((A & B) & C) & D))
                        reg_fstate <= state1;
                    else if ((((~(A) | ~(B)) | ~(C)) | ~(D)))
                        reg_fstate <= state0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state0;
                end
                state3: begin
                    reg_fstate <= state4;

                    CE <= 1'b1;
                end
                state1: begin
                    if (PBGNT)
                        reg_fstate <= state2;
                    else if (~(PBGNT))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    PBREQ <= 1'b1;
                end
                state2: begin
                    if (MACK)
                        reg_fstate <= state3;
                    else if (~(MACK))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    CMREQ <= 1'b1;

                    CNTLD <= 1'b1;
                end
                state4: begin
                    if (~(CONT))
                        reg_fstate <= state0;
                    else if (CONT)
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;
                end
                state5: begin
                    if (MACK)
                        reg_fstate <= state3;
                    else if (~(MACK))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;
                end
                default: begin
                    PBREQ <= 1'bx;
                    CMREQ <= 1'bx;
                    CE <= 1'bx;
                    CNTLD <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // HW3Q6
